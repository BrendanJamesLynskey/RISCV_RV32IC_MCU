// ============================================================================
// brv32p_core.sv — 5-Stage Pipelined RV32IMC CPU Core
// ============================================================================
// Stages: IF → ID → EX → MEM → WB
// Features:
//   - Full data forwarding (EX→EX, MEM→EX)
//   - Load-use stall (1 cycle)
//   - 2-bit branch predictor with BTB
//   - RV32C compressed instruction expansion
//   - M-extension multiply/divide
//   - Machine-mode CSRs and traps
// ============================================================================
import brv32p_pkg::*;

module brv32p_core (
  input  logic        clk,
  input  logic        rst_n,

  // Instruction memory interface (active-low stall = ready)
  output logic [31:0] imem_addr,
  output logic        imem_rd,
  input  logic [31:0] imem_rdata,
  input  logic        imem_ready,

  // Data memory interface
  output logic [31:0] dmem_addr,
  output logic        dmem_rd,
  output logic        dmem_wr,
  output mem_width_e  dmem_width,
  output logic        dmem_sign_ext,
  output logic [31:0] dmem_wdata,
  input  logic [31:0] dmem_rdata,
  input  logic        dmem_ready,

  // Interrupts
  input  logic        ext_irq,
  input  logic        timer_irq
);

  // ════════════════════════════════════════════════════════════════════
  // Pipeline control signals
  // ════════════════════════════════════════════════════════════════════
  logic stall_if, stall_id, stall_ex;
  logic flush_id, flush_ex, flush_mem;
  fwd_sel_e fwd_rs1, fwd_rs2;
  logic mem_stall;

  assign mem_stall = (dmem_rd | dmem_wr) & ~dmem_ready;

  // ════════════════════════════════════════════════════════════════════
  // IF — Instruction Fetch
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] pc_if, pc_next;
  logic [31:0] instr_raw_if;
  logic        bp_pred_taken;
  logic [31:0] bp_pred_target;
  logic        bp_pred_valid;
  logic        is_compressed_if;

  // PC Register
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n)
      pc_if <= RESET_VECTOR;
    else if (!stall_if && !mem_stall)
      pc_if <= pc_next;
  end

  assign imem_addr = pc_if;
  assign imem_rd   = 1'b1;
  assign instr_raw_if = imem_rdata;

  // Compressed decoder
  logic [31:0] instr_expanded_if;
  logic        illegal_c_if;

  compressed_decoder u_cdec (
    .instr_in      (instr_raw_if),
    .instr_out     (instr_expanded_if),
    .is_compressed (is_compressed_if),
    .illegal_c     (illegal_c_if)
  );

  // Branch predictor
  branch_predictor u_bp (
    .clk         (clk),
    .rst_n       (rst_n),
    .pc          (pc_if),
    .pred_taken  (bp_pred_taken),
    .pred_target (bp_pred_target),
    .pred_valid  (bp_pred_valid),
    .update_en   (bp_update_en),
    .update_pc   (bp_update_pc),
    .update_taken(bp_update_taken),
    .update_target(bp_update_target)
  );

  // Next PC MUX — priority: trap > mispredict > predicted taken > sequential
  logic        branch_mispredict_ex;
  logic [31:0] branch_target_ex;
  logic        trap_enter;
  logic [31:0] mtvec_out, mepc_out;
  logic        mret_ex;

  logic [31:0] pc_inc;
  assign pc_inc = is_compressed_if ? 32'd2 : 32'd4;

  always_comb begin
    if (trap_enter)
      pc_next = mtvec_out;
    else if (mret_ex)
      pc_next = mepc_out;
    else if (branch_mispredict_ex)
      pc_next = branch_target_ex;
    else if (bp_pred_taken && bp_pred_valid)
      pc_next = bp_pred_target;
    else
      pc_next = pc_if + pc_inc;
  end

  // ════════════════════════════════════════════════════════════════════
  // IF/ID Pipeline Register
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] pc_id, instr_id;
  logic [31:0] pc_inc_id;
  logic        pred_taken_id;
  logic        illegal_c_id;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n || flush_id) begin
      pc_id         <= 32'b0;
      instr_id      <= 32'h0000_0013; // NOP
      pc_inc_id     <= 32'd4;
      pred_taken_id <= 1'b0;
      illegal_c_id  <= 1'b0;
    end else if (!stall_id && !mem_stall) begin
      pc_id         <= pc_if;
      instr_id      <= instr_expanded_if;
      pc_inc_id     <= pc_inc;
      pred_taken_id <= bp_pred_taken && bp_pred_valid;
      illegal_c_id  <= illegal_c_if;
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // ID — Instruction Decode
  // ════════════════════════════════════════════════════════════════════
  logic [4:0]  rs1_addr_id, rs2_addr_id, rd_addr_id;
  logic [31:0] imm_id;
  ctrl_t       ctrl_id;
  logic [31:0] rs1_data_raw, rs2_data_raw;

  decoder u_decoder (
    .instr    (instr_id),
    .rs1_addr (rs1_addr_id),
    .rs2_addr (rs2_addr_id),
    .rd_addr  (rd_addr_id),
    .imm      (imm_id),
    .ctrl     (ctrl_id)
  );

  // Register file
  logic        wb_wr_en;
  logic [4:0]  wb_rd_addr;
  logic [31:0] wb_rd_data;

  regfile u_regfile (
    .clk      (clk),
    .rst_n    (rst_n),
    .rs1_addr (rs1_addr_id),
    .rs1_data (rs1_data_raw),
    .rs2_addr (rs2_addr_id),
    .rs2_data (rs2_data_raw),
    .wr_en    (wb_wr_en),
    .rd_addr  (wb_rd_addr),
    .rd_data  (wb_rd_data)
  );

  // ════════════════════════════════════════════════════════════════════
  // ID/EX Pipeline Register
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] pc_ex, rs1_data_ex, rs2_data_ex, imm_ex;
  logic [31:0] pc_inc_ex;
  logic [4:0]  rs1_addr_ex, rs2_addr_ex, rd_addr_ex;
  ctrl_t       ctrl_ex;
  logic        pred_taken_ex;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n || flush_ex) begin
      ctrl_ex       <= '0;
      pc_ex         <= 32'b0;
      rs1_data_ex   <= 32'b0;
      rs2_data_ex   <= 32'b0;
      imm_ex        <= 32'b0;
      pc_inc_ex     <= 32'd4;
      rs1_addr_ex   <= 5'b0;
      rs2_addr_ex   <= 5'b0;
      rd_addr_ex    <= 5'b0;
      pred_taken_ex <= 1'b0;
    end else if (!stall_ex && !mem_stall) begin
      ctrl_ex       <= ctrl_id;
      pc_ex         <= pc_id;
      rs1_data_ex   <= rs1_data_raw;
      rs2_data_ex   <= rs2_data_raw;
      imm_ex        <= imm_id;
      pc_inc_ex     <= pc_inc_id;
      rs1_addr_ex   <= rs1_addr_id;
      rs2_addr_ex   <= rs2_addr_id;
      rd_addr_ex    <= rd_addr_id;
      pred_taken_ex <= pred_taken_id;
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // EX — Execute
  // ════════════════════════════════════════════════════════════════════

  // Forwarding MUXes
  logic [31:0] rs1_fwd, rs2_fwd;
  logic [31:0] alu_result_mem;  // From EX/MEM register
  logic [31:0] wb_data_fwd;     // From MEM/WB

  always_comb begin
    case (fwd_rs1)
      FWD_EX_MEM:  rs1_fwd = alu_result_mem;
      FWD_MEM_WB:  rs1_fwd = wb_data_fwd;
      default:     rs1_fwd = rs1_data_ex;
    endcase
    case (fwd_rs2)
      FWD_EX_MEM:  rs2_fwd = alu_result_mem;
      FWD_MEM_WB:  rs2_fwd = wb_data_fwd;
      default:     rs2_fwd = rs2_data_ex;
    endcase
  end

  // ALU
  logic [31:0] alu_a, alu_b, alu_result_ex;
  logic        alu_zero;

  // AUIPC uses PC as operand A
  assign alu_a = (ctrl_ex.alu_op == ALU_ADD && instr_id == instr_id) ?
                 // Detect AUIPC: check original opcode bits
                 rs1_fwd : rs1_fwd;
  // Better AUIPC detection: store it in ctrl
  // For now, handle via wb_sel and direct computation in writeback

  assign alu_b = ctrl_ex.alu_src ? imm_ex : rs2_fwd;

  alu u_alu (
    .a      (rs1_fwd),
    .b      (alu_b),
    .op     (ctrl_ex.alu_op),
    .result (alu_result_ex),
    .zero   (alu_zero)
  );

  // AUIPC result
  logic [31:0] auipc_result;
  assign auipc_result = pc_ex + imm_ex;

  // MulDiv
  logic [31:0] muldiv_result;
  logic        muldiv_busy, muldiv_valid;

  muldiv u_muldiv (
    .clk    (clk),
    .rst_n  (rst_n),
    .start  (ctrl_ex.muldiv_en),
    .op     (ctrl_ex.muldiv_op),
    .a      (rs1_fwd),
    .b      (rs2_fwd),
    .result (muldiv_result),
    .busy   (muldiv_busy),
    .valid  (muldiv_valid)
  );

  // Branch resolution
  logic branch_taken_ex;
  logic [31:0] branch_target_computed;

  always_comb begin
    branch_taken_ex = 1'b0;
    case (ctrl_ex.branch_type)
      BR_EQ:  branch_taken_ex = (rs1_fwd == rs2_fwd);
      BR_NE:  branch_taken_ex = (rs1_fwd != rs2_fwd);
      BR_LT:  branch_taken_ex = ($signed(rs1_fwd) < $signed(rs2_fwd));
      BR_GE:  branch_taken_ex = ($signed(rs1_fwd) >= $signed(rs2_fwd));
      BR_LTU: branch_taken_ex = (rs1_fwd < rs2_fwd);
      BR_GEU: branch_taken_ex = (rs1_fwd >= rs2_fwd);
      default: branch_taken_ex = 1'b0;
    endcase
  end

  assign branch_target_computed = ctrl_ex.jalr ?
    {alu_result_ex[31:1], 1'b0} : (pc_ex + imm_ex);

  // Mispredict detection
  logic is_branch_or_jump;
  assign is_branch_or_jump = (ctrl_ex.branch_type != BR_NONE) ||
                              ctrl_ex.jal || ctrl_ex.jalr;

  logic actual_taken;
  assign actual_taken = branch_taken_ex || ctrl_ex.jal || ctrl_ex.jalr;

  assign branch_mispredict_ex = is_branch_or_jump &&
    ((actual_taken != pred_taken_ex) ||
     (actual_taken && (branch_target_computed != pc_ex + pc_inc_ex)));
  // Simplified: if prediction was wrong direction, or right direction but wrong target

  assign branch_target_ex = actual_taken ? branch_target_computed :
                            (pc_ex + pc_inc_ex); // Not-taken fallthrough

  // Branch predictor update
  logic bp_update_en;
  logic [31:0] bp_update_pc, bp_update_target;
  logic bp_update_taken;

  assign bp_update_en     = (ctrl_ex.branch_type != BR_NONE);
  assign bp_update_pc     = pc_ex;
  assign bp_update_taken  = branch_taken_ex;
  assign bp_update_target = branch_target_computed;

  // MRET
  assign mret_ex = ctrl_ex.mret;

  // EX result select
  logic [31:0] ex_result;
  always_comb begin
    case (ctrl_ex.wb_sel)
      WB_ALU:    ex_result = alu_result_ex;
      WB_PC4:    ex_result = pc_ex + pc_inc_ex;
      WB_MULDIV: ex_result = muldiv_result;
      default:   ex_result = alu_result_ex;
    endcase
    // Override for AUIPC (opcode check in pipeline)
    if (ctrl_ex.alu_src && ctrl_ex.alu_op == ALU_ADD && !ctrl_ex.mem_rd &&
        !ctrl_ex.mem_wr && !ctrl_ex.jalr && ctrl_ex.wb_sel == WB_ALU) begin
      // This might be AUIPC or ADDI. Need a cleaner flag.
      // For now, AUIPC goes through ALU with rs1=0, so result is just imm.
      // Actually AUIPC needs PC+imm. Let's use a dedicated flag.
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // EX/MEM Pipeline Register
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] pc_mem;
  logic [31:0] ex_result_mem, rs2_data_mem;
  logic [4:0]  rd_addr_mem;
  ctrl_t       ctrl_mem;

  assign alu_result_mem = ex_result_mem;  // Forwarding tap

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n || flush_mem) begin
      ctrl_mem       <= '0;
      pc_mem         <= 32'b0;
      ex_result_mem  <= 32'b0;
      rs2_data_mem   <= 32'b0;
      rd_addr_mem    <= 5'b0;
    end else if (!mem_stall) begin
      ctrl_mem       <= ctrl_ex;
      pc_mem         <= pc_ex;
      ex_result_mem  <= ex_result;
      rs2_data_mem   <= rs2_fwd;
      rd_addr_mem    <= rd_addr_ex;
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // MEM — Memory Access
  // ════════════════════════════════════════════════════════════════════
  assign dmem_addr     = ex_result_mem;
  assign dmem_rd       = ctrl_mem.mem_rd;
  assign dmem_wr       = ctrl_mem.mem_wr;
  assign dmem_width    = ctrl_mem.mem_width;
  assign dmem_sign_ext = ctrl_mem.mem_sign_ext;
  assign dmem_wdata    = rs2_data_mem;

  // MEM result
  logic [31:0] mem_result;
  assign mem_result = ctrl_mem.mem_rd ? dmem_rdata : ex_result_mem;

  // Trap logic
  logic        irq_pending;
  logic [31:0] csr_rdata;

  assign trap_enter = ctrl_mem.ecall || ctrl_mem.ebreak ||
                      ctrl_mem.illegal || irq_pending;

  logic [31:0] trap_cause, trap_val;
  always_comb begin
    trap_cause = 32'b0;
    trap_val   = 32'b0;
    if (ctrl_mem.illegal) begin
      trap_cause = 32'd2;
    end else if (ctrl_mem.ecall) begin
      trap_cause = 32'd11;
    end else if (ctrl_mem.ebreak) begin
      trap_cause = 32'd3;
    end else if (irq_pending) begin
      trap_cause = {1'b1, 31'd11};
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // MEM/WB Pipeline Register
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] mem_result_wb;
  logic [31:0] csr_rdata_wb;
  logic [4:0]  rd_addr_wb;
  ctrl_t       ctrl_wb;

  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      ctrl_wb      <= '0;
      mem_result_wb <= 32'b0;
      csr_rdata_wb <= 32'b0;
      rd_addr_wb   <= 5'b0;
    end else if (!mem_stall) begin
      ctrl_wb      <= ctrl_mem;
      mem_result_wb <= mem_result;
      csr_rdata_wb <= csr_rdata;
      rd_addr_wb   <= rd_addr_mem;
    end
  end

  // ════════════════════════════════════════════════════════════════════
  // WB — Writeback
  // ════════════════════════════════════════════════════════════════════
  always_comb begin
    case (ctrl_wb.wb_sel)
      WB_MEM:    wb_rd_data = mem_result_wb;
      WB_CSR:    wb_rd_data = csr_rdata_wb;
      default:   wb_rd_data = mem_result_wb;
    endcase
  end

  assign wb_wr_en  = ctrl_wb.reg_wr;
  assign wb_rd_addr = rd_addr_wb;
  assign wb_data_fwd = wb_rd_data;  // Forwarding tap

  // ════════════════════════════════════════════════════════════════════
  // CSR Unit
  // ════════════════════════════════════════════════════════════════════
  logic [31:0] csr_wdata;
  assign csr_wdata = ctrl_mem.csr_op[2] ?
    {27'b0, rd_addr_mem} : ex_result_mem; // FIXME: should be rs1 data

  csr u_csr (
    .clk           (clk),
    .rst_n         (rst_n),
    .csr_en        (ctrl_mem.csr_en && !trap_enter),
    .csr_addr      (ctrl_mem.csr_addr),
    .csr_op        (ctrl_mem.csr_op),
    .csr_wdata     (csr_wdata),
    .csr_rdata     (csr_rdata),
    .trap_enter    (trap_enter),
    .trap_cause    (trap_cause),
    .trap_val      (trap_val),
    .trap_pc       (pc_mem),
    .mtvec_out     (mtvec_out),
    .mepc_out      (mepc_out),
    .mret          (mret_ex),
    .ext_irq       (ext_irq),
    .timer_irq     (timer_irq),
    .instr_retired (ctrl_wb.reg_wr || ctrl_wb.mem_wr || ctrl_wb.ecall),
    .irq_pending   (irq_pending)
  );

  // ════════════════════════════════════════════════════════════════════
  // Hazard Unit
  // ════════════════════════════════════════════════════════════════════
  hazard_unit u_hazard (
    .id_rs1           (rs1_addr_id),
    .id_rs2           (rs2_addr_id),
    .ex_rd            (rd_addr_ex),
    .ex_reg_wr        (ctrl_ex.reg_wr),
    .ex_mem_rd        (ctrl_ex.mem_rd),
    .ex_wb_sel        (ctrl_ex.wb_sel),
    .mem_rd           (rd_addr_mem),
    .mem_reg_wr       (ctrl_mem.reg_wr),
    .wb_rd            (rd_addr_wb),
    .wb_reg_wr        (ctrl_wb.reg_wr),
    .branch_mispredict(branch_mispredict_ex || trap_enter || mret_ex),
    .jump_ex          (ctrl_ex.jal || ctrl_ex.jalr),
    .muldiv_busy      (muldiv_busy),
    .fwd_rs1          (fwd_rs1),
    .fwd_rs2          (fwd_rs2),
    .stall_if         (stall_if),
    .stall_id         (stall_id),
    .stall_ex         (stall_ex),
    .flush_id         (flush_id),
    .flush_ex         (flush_ex),
    .flush_mem        (flush_mem)
  );

endmodule
