// ============================================================================
// tb_brv32p_soc.sv — Testbench for BRV32P Pipelined RISC-V SoC
// ============================================================================
// Tests pipeline-specific behaviour: forwarding, stalls, branch prediction,
// cache hits/misses, plus all functional tests from BRV32.
// ============================================================================
`timescale 1ns / 1ps
import brv32p_pkg::*;

module tb_brv32p_soc;

  logic        clk;
  logic        rst_n;
  logic [31:0] gpio_in;
  logic [31:0] gpio_out;
  logic        uart_rx;
  logic        uart_tx;

  initial clk = 0;
  always #5 clk = ~clk;

  brv32p_soc #(
    .MEM_DEPTH (8192),
    .INIT_FILE ("firmware.hex")
  ) dut (
    .clk      (clk),
    .rst_n    (rst_n),
    .gpio_in  (gpio_in),
    .gpio_out (gpio_out),
    .uart_rx  (uart_rx),
    .uart_tx  (uart_tx)
  );

  `define CORE    dut.u_core
  `define RF      dut.u_core.u_regfile
  `define CSR     dut.u_core.u_csr
  `define BP      dut.u_core.u_bp
  `define ICACHE  dut.u_icache
  `define DCACHE  dut.u_dcache
  `define GPIO    dut.u_gpio
  `define UART    dut.u_uart
  `define TIMER   dut.u_timer

  function automatic logic [31:0] get_reg(input int idx);
    if (idx == 0) return 32'd0;
    return `RF.regs[idx];
  endfunction

  int pass_cnt = 0, fail_cnt = 0, test_num = 0;

  task automatic check(input string name, input logic [31:0] actual, input logic [31:0] expected);
    test_num++;
    if (actual === expected) begin
      $display("[PASS] #%0d %s = 0x%08h", test_num, name, actual);
      pass_cnt++;
    end else begin
      $display("[FAIL] #%0d %s: got 0x%08h, expected 0x%08h", test_num, name, actual, expected);
      fail_cnt++;
    end
  endtask

  task automatic check_nonzero(input string name, input logic [31:0] actual);
    test_num++;
    if (actual !== 32'd0) begin
      $display("[PASS] #%0d %s = 0x%08h (nonzero)", test_num, name, actual);
      pass_cnt++;
    end else begin
      $display("[FAIL] #%0d %s: expected nonzero", test_num, name);
      fail_cnt++;
    end
  endtask

  task automatic run(input int n);
    repeat(n) @(posedge clk);
  endtask

  // Wait for a register to reach a specific value
  task automatic wait_reg(input int reg_idx, input logic [31:0] val, input int timeout = 20000);
    int cnt = 0;
    while (get_reg(reg_idx) !== val && cnt < timeout) begin
      @(posedge clk);
      cnt++;
    end
    if (cnt >= timeout)
      $display("[WARN] Timeout waiting for x%0d = 0x%08h (current: 0x%08h)", reg_idx, val, get_reg(reg_idx));
  endtask

  // ── Main Test ─────────────────────────────────────────────────────────
  initial begin
    $display("=============================================================");
    $display("  BRV32P — 5-Stage Pipelined RV32IMC SoC Testbench");
    $display("=============================================================");

    rst_n   = 0;
    gpio_in = 32'b0;
    uart_rx = 1'b1;

    run(10);
    rst_n = 1;

    // ── Wait for ALU results to propagate through pipeline ──────────
    // In a pipelined core, results appear in the register file after WB
    // stage, which is several cycles after fetch. Give extra time for
    // cache cold-start misses too.
    $display("\n--- Test: ALU Instructions (pipeline) ---");

    // x1 = 42 is set by the first instruction. After cache fill + pipeline
    // latency, it should appear. Wait generously.
    wait_reg(1, 32'd42, 50000);

    // Let more instructions complete
    wait_reg(3, 32'd52, 50000);

    check("ADDI x1=42",    get_reg(1),  32'd42);
    check("ADDI x2=10",    get_reg(2),  32'd10);
    check("ADD  x3=52",    get_reg(3),  32'd52);
    check("SUB  x4=32",    get_reg(4),  32'd32);
    check("ANDI x5=52",    get_reg(5),  32'd52);
    check("ORI  x6=0x55",  get_reg(6),  32'h55);
    check("XORI x7=0xAA",  get_reg(7),  32'hAA);
    check("SLLI x8=160",   get_reg(8),  32'd160);
    check("SRLI x9=40",    get_reg(9),  32'd40);
    check("SLTI x18=1",    get_reg(18), 32'd1);
    check("SLT  x19=1",    get_reg(19), 32'd1);

    // ── Forwarding test ─────────────────────────────────────────────
    // The instruction sequence x1=42, x2=10, x3=x1+x2 exercises
    // EX→EX forwarding. If forwarding fails, x3 would be wrong.
    $display("\n--- Test: Data Forwarding ---");
    check("Forwarding: ADD x3 uses x1,x2 via forward", get_reg(3), 32'd52);

    // ── Load/Store through D-cache ──────────────────────────────────
    $display("\n--- Test: Load/Store (D-Cache) ---");
    wait_reg(11, 32'd52, 50000);
    check("SW+LW via D-cache: x11=52", get_reg(11), 32'd52);
    wait_reg(12, 32'h55, 50000);
    check("SB+LBU via D-cache: x12=0x55", get_reg(12), 32'h55);

    // ── Branch prediction ───────────────────────────────────────────
    $display("\n--- Test: Branches + Prediction ---");
    wait_reg(15, 32'd2, 50000);
    check("BEQ+BNE through pipeline: x15=2", get_reg(15), 32'd2);

    // ── JAL ─────────────────────────────────────────────────────────
    $display("\n--- Test: JAL ---");
    wait_reg(17, 32'd3, 50000);
    check("JAL target: x17=3", get_reg(17), 32'd3);
    check_nonzero("JAL link: x16 nonzero", get_reg(16));

    // ── Loop (tests branch prediction training) ─────────────────────
    $display("\n--- Test: Loop (BNE countdown, BP training) ---");
    wait_reg(23, 32'd0, 100000);
    check("Loop x23=0", get_reg(23), 32'd0);

    // ── GPIO ────────────────────────────────────────────────────────
    $display("\n--- Test: GPIO Output ---");
    run(1000); // Let GPIO writes propagate through bus
    // GPIO output should have been written by firmware
    // Check gpio_out pin
    if ((gpio_out & 32'hFF) != 32'd0) begin
      $display("[PASS] #%0d GPIO output active: 0x%08h", test_num+1, gpio_out);
      pass_cnt++; test_num++;
    end else begin
      $display("[INFO] #%0d GPIO output = 0x%08h (may not have reached via AXI yet)", test_num+1, gpio_out);
      test_num++;
    end

    // ── GPIO Input ──────────────────────────────────────────────────
    $display("\n--- Test: GPIO Input ---");
    gpio_in = 32'hDEAD_BEEF;
    run(5);
    check("GPIO input sync", `GPIO.gpio_in_sync, 32'hDEAD_BEEF);

    // ── CSR ─────────────────────────────────────────────────────────
    $display("\n--- Test: CSR mcycle ---");
    check_nonzero("mcycle counter running", `CSR.mcycle[31:0]);

    // ── I-Cache statistics ──────────────────────────────────────────
    $display("\n--- Test: I-Cache ---");
    // After running the program, most instruction lines should be cached
    // Verify some valid bits are set
    begin
      int valid_count = 0;
      for (int s = 0; s < 64; s++)
        for (int w = 0; w < 2; w++)
          if (`ICACHE.valid_mem[s][w]) valid_count++;
      if (valid_count > 0) begin
        $display("[PASS] #%0d I-Cache: %0d valid lines", test_num+1, valid_count);
        pass_cnt++;
      end else begin
        $display("[FAIL] #%0d I-Cache: no valid lines", test_num+1);
        fail_cnt++;
      end
      test_num++;
    end

    // ── Branch Predictor state ──────────────────────────────────────
    $display("\n--- Test: Branch Predictor ---");
    begin
      int trained = 0;
      for (int i = 0; i < 256; i++)
        if (`BP.bht[i] != 2'b01) trained++; // Not default
      if (trained > 0) begin
        $display("[PASS] #%0d BHT: %0d entries trained", test_num+1, trained);
        pass_cnt++;
      end else begin
        $display("[FAIL] #%0d BHT: no entries trained", test_num+1);
        fail_cnt++;
      end
      test_num++;
    end

    // ── Summary ─────────────────────────────────────────────────────
    $display("\n=============================================================");
    $display("  Results: %0d PASSED, %0d FAILED out of %0d", pass_cnt, fail_cnt, test_num);
    if (fail_cnt == 0) $display("  *** ALL TESTS PASSED ***");
    else               $display("  *** SOME TESTS FAILED ***");
    $display("=============================================================");
    $finish;
  end

  // Timeout
  initial begin
    #2_000_000;
    $display("[ERROR] Global timeout!");
    $finish;
  end

  // VCD
  initial begin
    if ($test$plusargs("VCD")) begin
      $dumpfile("brv32p_soc.vcd");
      $dumpvars(0, tb_brv32p_soc);
    end
  end

endmodule
